`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:25:22 11/03/2024 
// Design Name: 
// Module Name:    ANGLE_CALCULATOR 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ANGLE_CALCULATOR(
    input [2:0] rt,
    input [2:0] rd,
    input [2:0] ld,
    input [2:0] lt,
    input [2:0] gx,
    input [2:0] gy,
    input xDir,
    input yDir
    );


endmodule
